--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
--                                                                            --
-- top heading: TM FAST Library package                                       --
--                                                                            --
-- filename:    TFL_FAST_USER_LIB_p.vhd                                       --
--                                                                            --                                                           
-- revision:    see TFL_FAST_USER_LIB_LOG_VER_CC                              --
--                                                                            --
-- copyright:   Siemens AG, Digital Industries, Factory Automation            --
--                                                                            --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


package TFL_FAST_USER_LIB_p is


  -- logic version
  constant  TFL_FAST_USER_LIB_LOG_VER_CC:  string ( 1 to 9 ) := "V03.00.00"; -- TFL logic-version format: <TYPE>xx.yy.zz

end package TFL_FAST_USER_LIB_p;
